module fifo_goertzel_tb();











endmodule