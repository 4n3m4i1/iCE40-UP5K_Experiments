

module top 
(
    input       button,
    output wire LED
);


/*
module SR_DB
#(
    parameter SYSCLK_FREQ = 24000000,
    parameter DEBOUNCE_DELAY = 0.150
)(
    input       clk,
    input       D,
    output reg  Q
);
*/

endmodule